module datapath
(
	input		USER_CLK,
	input		
